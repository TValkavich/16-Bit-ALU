`timescale 1ns/1ns //timescale of 1 nanosecond

module testBench(); //calls to test my ALU
	wire[15:0] A, B, Set, F, Cout;
	wire Sub, Op1, Op2, Less, Cin;
	testALU16 test (F, Cout, Set, Less, A, B, Cin, Sub, Op1, Op2);
	ALU16 alu (F, Cout, Set, Less, A, B, Cin, Sub, Op1, Op2);
endmodule

module testALU16(F, Cout, Set, Less, A, B, Cin, Sub, Op1, Op2); //inputs values into 16-bit ALU
	input [15:0] F, Set, Cout;
	output [15:0] A, B;
	output Cin, Sub, Op1, Op2, Less;
	reg [15:0] A, B;
	reg Cin, Sub, Op1, Op2, Less;    
	initial
		begin
			$monitor($time, ,"A=%d, B=%d, Cin=%b, F=%d, Cout=%b, Set=%b, Sub=%b, Op1=%b, Op2=%b, Less=%b", A, B, Cin,F, Cout, Set, Sub, Op1, Op2, Less);
			$display($time, ,"A=%d, B=%d, Cin=%b, F=%d, Cout=%b, Set=%b, Sub=%b, Op1=%b, Op2=%b, Less=%b", A, B, Cin,F, Cout, Set, Sub, Op1, Op2, Less);
			
			//1000 RANDOM INPUTS BELOW

			//AND - Postive and Neagtive Inputs with a 100 nanosecond delay
			#100 A =4555; B =1; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1; B =1; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =637; B =120; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3555; B =1245; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =21982; B =4750; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =50; B =-20; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2345; B =7303; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =26; B =2685; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =864; B =8231; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =245; B =5160; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8975; B =0789; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =124; B =6483; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3; B =3385; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =684; B =5873; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =346; B =7120; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =895; B =5193; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =246; B =3476; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =908; B =2849; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7654; B =2430; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1245; B =5642; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =688; B =7777; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =674; B =9926; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =365; B =7687; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =376; B =9850; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =745; B =2603; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2324; B =2899; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1235; B =7217; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =677; B =0202; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5; B =1478; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =54; B =9925; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =34; B =2882; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =876; B =9119; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =12; B =2121; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1; B =2294; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =786; B =7178; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8; B =7697; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6; B =7745; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =57; B =6641; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =12; B =4907; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4356; B =8390; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =43; B =0487; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =764; B =5912; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =467; B =5505; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2345; B =0193; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =78; B =8625; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =287; B =6860; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =798; B =7484; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =34; B =3002; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =65; B =4151; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =687; B =3534; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =76; B =7232; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =234; B =2393; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =345; B =5207; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =56; B =1630; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =546; B =8433; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =345; B =2113; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =76; B =7843; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1; B =8587; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7; B =4995; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5; B =9706; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4; B =5790; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =234; B =0381; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =765; B =2540; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7666; B =8524; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =222; B =0979; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =222; B =7151; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =111; B =3598; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =222; B =7050; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =457; B =4569; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =654; B =1903; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7446; B =0089; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =676; B =8629; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =543; B =3808; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =676; B =5188; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =567; B =8503; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =567; B =5580; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =876; B =4349; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8765; B =1479; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =345; B =5069; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =454; B =3081; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4356; B =1663; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =452; B =2997; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =123; B =1841; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =767; B =0412; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =654; B =8692; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =67; B =0249; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =98; B =8818; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3; B =6096; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =376; B =3109; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =87; B =8537; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =124; B =4848; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =45; B =8458; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =67; B =4009; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =87; B =7565; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =13; B =1359; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =12; B =1553; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =346; B =9115; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =67; B =3430; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =654; B =4652; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =675; B =9382; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =12; B =9266; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =346; B =9542; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =658; B =1122; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =876; B =4836; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =124; B =7455; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3257; B =0144; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =765; B =0884; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =698; B =9920; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =12; B =8582; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =77; B =4202; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =876; B =2973; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4356; B =6009; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =987; B =3737; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =54; B =0189; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =436; B =6862; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =765; B =1395; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =98; B =3633; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =908; B =6355; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =865; B =6497; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =658; B =6453; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =234; B =1267; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =357; B =8536; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =797; B =8364; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =124; B =9890; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5; B =2134; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =45; B =8755; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =12; B =0463; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =87; B =3654; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =543; B =4793; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7; B =0101; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8765; B =2961; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6543; B =3308; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =35; B =5526; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =56; B =2910; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =768; B =0109; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5643; B =1426; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =43; B =4198; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =567; B =4676; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =765; B =3185; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =543; B =1075; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =436; B =9216; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =765; B =9574; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1; B =6854; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =234; B =4709; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =56; B =2419; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =543; B =8938; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =568; B =2524; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =344; B =7207; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6544; B =8359; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1111; B =5389; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5876; B =3457; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6543; B =4052; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =543; B =3231; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =657; B =8911; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =67; B =7184; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =890; B =6382; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =40; B =0464; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4345; B =2146; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =679; B =3363; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9876; B =7832; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =432; B =4885; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =347; B =5696; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6798; B =6689; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =876; B =4079; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =640; B =1918; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8765; B =7354; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =543; B =5104; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =12; B =7065; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =123; B =8727; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2; B =5429; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7; B =6311; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =900; B =3079; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7654; B =2005; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =453; B =8947; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =43; B =4443; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =457; B =9315; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =67; B =5682; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5; B =1360; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8; B =4432; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =98; B =8700; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7654; B =4680; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =32; B =1275; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =84; B =9577; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =723; B =5051; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =43; B =5506; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =458; B =5849; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =908; B =6181; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			#100 A =65; B =1870; Sub = 0;Op1 = 0; Op2 = 0; Cin = 0; Less = 0;
			
			//OR - Postive and Neagtive Inputs with a 100 nanosecond delay
			#100 A =6718; B =1; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1; B =1; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =637; B =120; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3555; B =1245; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =21982; B =4750; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =50; B =-20; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7546; B =3839; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2267; B =1911; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9186; B =8119; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0029; B =9879; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5892; B =0124; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2803; B =6042; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1463; B =0654; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2125; B =8259; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9593; B =1905; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0803; B =7727; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7345; B =7317; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5036; B =1527; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4008; B =6228; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5908; B =2183; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2413; B =7344; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9284; B =6768; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8840; B =0552; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0064; B =0645; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7109; B =1476; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6945; B =4920; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7889; B =4855; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5413; B =8953; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2047; B =9493; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4208; B =6639; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9860; B =8241; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9191; B =7418; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2250; B =6215; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3915; B =8339; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2502; B =6050; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3256; B =9287; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0774; B =6565; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6826; B =4253; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0181; B =3448; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3669; B =3204; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4858; B =8738; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3068; B =0784; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7856; B =6271; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1729; B =2793; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7956; B =2445; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5733; B =7767; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9054; B =0025; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3164; B =3732; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5267; B =1821; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6460; B =7206; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3673; B =2116; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6108; B =3457; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7820; B =3485; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3111; B =9041; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9934; B =6244; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1049; B =9478; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1380; B =5432; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0048; B =3613; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7951; B =9896; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1840; B =1543; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3004; B =6827; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5448; B =7258; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0288; B =8165; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3787; B =5084; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8252; B =7867; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4167; B =7236; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0568; B =3780; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2713; B =8671; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1981; B =4584; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7530; B =4554; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0590; B =5238; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5284; B =4048; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5313; B =1048; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8267; B =5948; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2950; B =0380; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6754; B =6493; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0897; B =9308; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9907; B =8789; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8198; B =4820; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1706; B =6105; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8353; B =7895; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6904; B =0236; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3304; B =0949; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9556; B =1136; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0395; B =2903; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1016; B =3418; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9043; B =6345; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8444; B =7267; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1432; B =9239; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9909; B =7070; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7027; B =8123; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4064; B =1880; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5432; B =9822; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6195; B =8278; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6123; B =7256; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0861; B =8550; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0668; B =7126; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2793; B =4790; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6806; B =4866; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8180; B =1531; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9068; B =3593; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7707; B =3387; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8375; B =3998; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6804; B =6179; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7046; B =9594; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9826; B =1526; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2859; B =1641; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1619; B =8536; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6281; B =2615; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0131; B =2950; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5013; B =4435; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1298; B =2636; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3636; B =9171; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6819; B =5063; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5124; B =1365; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1065; B =0967; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7517; B =2445; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6411; B =2617; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0894; B =3273; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2506; B =6042; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0165; B =8203; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5259; B =6139; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0711; B =3837; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6447; B =1961; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4537; B =4798; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2755; B =8537; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0431; B =3959; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1451; B =9069; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3691; B =6545; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2714; B =6112; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4906; B =0103; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5670; B =2230; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0154; B =6160; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5590; B =0051; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0007; B =5675; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8859; B =9081; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0488; B =8851; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4721; B =7994; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7946; B =9750; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0179; B =1228; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7017; B =6277; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3142; B =6335; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2907; B =1733; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8360; B =7872; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7951; B =1915; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7523; B =9992; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4513; B =3810; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7847; B =1615; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0137; B =6025; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7356; B =1752; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4641; B =1572; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7156; B =1326; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0547; B =9245; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1231; B =7605; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8173; B =6910; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5735; B =9936; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0832; B =2792; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0738; B =8222; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7095; B =2612; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0767; B =3845; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2083; B =3467; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2495; B =0415; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2254; B =2719; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4666; B =1409; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5451; B =1394; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4194; B =9488; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3009; B =0625; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8325; B =7786; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4775; B =6106; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7236; B =9350; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1133; B =3133; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0794; B =4874; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7707; B =4228; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3296; B =9353; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1815; B =0767; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3949; B =7951; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2223; B =3124; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1311; B =8536; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4453; B =7049; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0633; B =4385; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5575; B =3813; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7690; B =5135; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7117; B =2967; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5615; B =0593; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3852; B =6189; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2318; B =9660; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5936; B =5907; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0350; B =7183; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0073; B =3573; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1161; B =8725; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0828; B =6098; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1071; B =0092; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4869; B =0526; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4431; B =5109; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9907; B =9800; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4156; B =6863; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =822; B =004; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =626; B =453; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =011; B =348; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =369; B =304; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =488; B =838; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =368; B =084; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =756; B =621; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =129; B =793; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =756; B =245; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =533; B =767; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			#100 A =904; B =025; Sub = 0;Op1 = 0; Op2 = 1; Cin = 0; Less = 0;
			
			//ADD - Postive and Neagtive Inputs with a 100 nanosecond delay
			#100 A =9631; B =1; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1; B =1; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =637; B =120; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3555; B =1245; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =21982; B =4750; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =50; B =-20; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6236; B =9897; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9966; B =5448; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1568; B =6231; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2431; B =1440; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9831; B =2953; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8723; B =1230; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4003; B =1737; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0149; B =9025; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6910; B =1924; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7902; B =6298; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0225; B =8711; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3917; B =8189; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7053; B =3122; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9942; B =9228; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2950; B =4922; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4157; B =2290; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4728; B =5396; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6122; B =0109; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5112; B =5520; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9554; B =4179; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5433; B =4229; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9215; B =3504; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0960; B =5146; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4566; B =0908; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6420; B =0932; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1179; B =9357; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2913; B =1251; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1044; B =3189; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2320; B =8347; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9132; B =0076; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2063; B =0112; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5375; B =4100; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9192; B =3905; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5618; B =2514; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7644; B =1818; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3129; B =7733; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7810; B =5086; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6788; B =6961; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6520; B =2511; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9486; B =4176; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1184; B =9292; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2010; B =6093; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3944; B =5588; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0041; B =8014; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1708; B =0991; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8194; B =7278; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6868; B =9388; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1050; B =7969; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2808; B =5009; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2524; B =1125; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5572; B =3145; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7269; B =7756; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3711; B =5580; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8722; B =9029; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8714; B =5409; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5475; B =7824; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6256; B =1969; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9939; B =9921; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1880; B =7940; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5299; B =9593; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2749; B =4329; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5477; B =3278; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6185; B =1553; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3894; B =6028; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9731; B =5447; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1952; B =7520; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0809; B =4378; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9408; B =5641; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0792; B =0441; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9104; B =8608; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1416; B =1585; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4774; B =0465; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8372; B =6827; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1775; B =3500; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0331; B =8503; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0251; B =6495; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0765; B =5650; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7496; B =4086; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6396; B =0934; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9523; B =4078; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4272; B =3519; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3295; B =6596; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4557; B =3745; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2968; B =2832; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4843; B =6136; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7222; B =2048; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9945; B =4619; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6660; B =2813; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7241; B =7732; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0639; B =3133; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2910; B =6206; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8551; B =8984; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3737; B =9570; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2938; B =9296; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4787; B =7372; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4189; B =3727; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4776; B =1290; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2093; B =8781; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0058; B =3291; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7336; B =8167; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1156; B =5183; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5619; B =4738; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2631; B =0961; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7035; B =3248; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0870; B =0079; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5365; B =9457; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3928; B =2112; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4084; B =2919; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8924; B =2341; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5831; B =7702; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7184; B =2978; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7908; B =0782; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8431; B =4201; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4446; B =2358; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9911; B =0423; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5014; B =2931; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3414; B =5748; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9183; B =8426; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5775; B =7370; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9722; B =9888; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1897; B =0585; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0042; B =7496; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4508; B =9642; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2546; B =1380; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0532; B =2505; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2523; B =1063; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6061; B =0089; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0468; B =7739; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7166; B =6260; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9793; B =9514; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7358; B =2508; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6786; B =5400; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8629; B =3896; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8526; B =2427; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6508; B =7947; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7788; B =2314; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4536; B =1526; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4379; B =9909; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7159; B =0154; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6638; B =7949; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5104; B =6384; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2752; B =6595; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0578; B =0032; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6047; B =6974; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7991; B =0041; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1103; B =9530; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7627; B =3496; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4586; B =4676; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1593; B =0786; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8195; B =8208; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2146; B =2658; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4239; B =6943; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7535; B =4316; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8167; B =2527; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7979; B =3793; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4405; B =4731; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8835; B =7020; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3150; B =4820; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0812; B =2907; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6456; B =0946; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8948; B =7423; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9285; B =8116; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6084; B =7157; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5364; B =5130; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7842; B =0841; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6769; B =9973; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4394; B =2977; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5132; B =8588; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5357; B =7767; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1903; B =7432; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7614; B =8268; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7628; B =8926; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5910; B =1085; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6141; B =7716; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2726; B =9102; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8464; B =6264; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8171; B =8150; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7172; B =7073; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9151; B =7308; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4676; B =7473; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7146; B =7473; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7449; B =8593; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3818; B =4918; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8894; B =7857; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5717; B =0579; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5714; B =7553; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6087; B =4161; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5816; B =3856; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5251; B =8987; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1889; B =8304; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3138; B =5343; Sub = 0;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			
			//SUB - Postive and Neagtive Inputs with a 100 nanosecond delay
			#100 A =7937; B =1; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1; B =1; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =637; B =120; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3555; B =1245; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =21982; B =4750; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =50; B =-20; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3665; B =0466; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7486; B =6942; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3410; B =1680; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6004; B =2988; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6542; B =5379; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4682; B =9930; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0546; B =8326; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2744; B =9082; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9327; B =1116; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9781; B =1576; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2210; B =4592; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2299; B =7459; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4654; B =3755; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5590; B =5593; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9208; B =8737; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2976; B =5529; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0007; B =7048; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8535; B =3242; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7508; B =0024; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3252; B =7827; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4031; B =5312; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8846; B =7003; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5683; B =1322; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9231; B =9086; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2675; B =9276; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9883; B =6156; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9773; B =5070; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0788; B =1133; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7503; B =1506; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9879; B =5254; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0927; B =8938; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7519; B =4312; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9930; B =1163; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5945; B =6320; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3208; B =5425; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7681; B =5503; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7645; B =5057; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4189; B =8685; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5119; B =4234; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6166; B =9442; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0634; B =6792; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7950; B =8228; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9578; B =9746; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3902; B =4108; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0541; B =8441; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7165; B =3256; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2288; B =8617; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4167; B =6426; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1092; B =2861; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6751; B =8393; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4851; B =2504; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7489; B =8405; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5991; B =9314; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3443; B =8794; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5716; B =6115; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9466; B =8347; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9584; B =3797; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0422; B =0692; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0584; B =9711; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5080; B =3065; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5364; B =1008; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9955; B =1700; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2121; B =3129; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1652; B =1085; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7479; B =2462; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9846; B =8632; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8865; B =7270; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8053; B =9960; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2565; B =9369; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4805; B =3721; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2025; B =9825; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3657; B =9416; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6832; B =3464; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9577; B =6308; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4813; B =7357; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0154; B =3952; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0101; B =3036; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0793; B =0687; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3988; B =9300; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1673; B =4237; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0114; B =5985; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5343; B =7497; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9315; B =3953; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2563; B =3367; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5486; B =3389; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1207; B =6005; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7997; B =2916; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9419; B =3049; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8087; B =1826; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2975; B =7253; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2169; B =3336; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4410; B =5683; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7212; B =0371; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1858; B =0577; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5143; B =2367; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2700; B =2861; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1390; B =0727; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2487; B =6464; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7553; B =6434; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4892; B =3364; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1759; B =6035; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4160; B =4061; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0290; B =0248; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5668; B =5067; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0728; B =7324; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9368; B =4640; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3400; B =1780; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9245; B =0101; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3729; B =2813; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6526; B =7050; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0174; B =9470; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7113; B =6063; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9785; B =7439; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4510; B =4445; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6839; B =6516; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4492; B =6014; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0605; B =1740; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1746; B =7064; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6838; B =3029; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6758; B =4124; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9300; B =9269; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5286; B =8328; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2118; B =6146; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0446; B =6626; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1152; B =5519; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2881; B =0912; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8442; B =3180; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3033; B =5616; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8718; B =0420; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9047; B =4164; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3354; B =3672; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3166; B =1340; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3218; B =9141; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7546; B =8999; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4611; B =4490; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1683; B =9907; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0459; B =7142; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3745; B =0792; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3189; B =7801; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5349; B =7172; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7541; B =4207; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4036; B =9061; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2686; B =3392; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4185; B =0722; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1230; B =9811; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8563; B =5650; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5647; B =1954; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3040; B =4585; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8385; B =1206; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5020; B =2303; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5664; B =8774; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2054; B =4504; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6407; B =8183; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1647; B =8618; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2765; B =1152; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8150; B =4153; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4776; B =6272; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2973; B =6675; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8980; B =6490; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4704; B =4972; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5260; B =1528; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4589; B =4423; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7572; B =6581; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4251; B =1890; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5449; B =1612; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2998; B =8220; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6795; B =8091; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8003; B =9281; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0424; B =3859; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =5252; B =3497; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6838; B =6294; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0221; B =3267; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1754; B =4158; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9330; B =6492; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =9833; B =1069; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2455; B =0815; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2013; B =1764; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2462; B =7024; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1551; B =0775; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2360; B =7315; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2865; B =2461; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0981; B =8153; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =6791; B =7871; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =4534; B =3599; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =8546; B =6452; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1726; B =6152; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =3430; B =5714; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =0628; B =0672; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =7517; B =8508; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =2876; B =8938; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			#100 A =1383; B =8859; Sub = 1;Op1 = 1; Op2 = 0; Cin = 0; Less = 0;
			
			//SLT - Postive and Neagtive Inputs with a 100 nanosecond delay
			#100 A =8264; B =1; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1; B =1; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =637; B =120; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3555; B =1245; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =21982; B =4750; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =50; B =-20; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =-50; B =-20; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0643; B =7939; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9694; B =4542; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9611; B =7708; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2233; B =8217; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9242; B =5519; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5822; B =3815; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1509; B =2547; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2634; B =9026; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4294; B =9202; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4976; B =0659; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4092; B =6178; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5797; B =2299; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4280; B =7243; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2060; B =2756; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4596; B =8695; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4542; B =7893; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0227; B =5146; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3702; B =3188; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9333; B =0181; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3753; B =0929; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7339; B =8386; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3883; B =2469; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6781; B =0019; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8135; B =8517; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3244; B =9865; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7571; B =2441; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8118; B =7793; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5425; B =5467; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4813; B =7873; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1420; B =8829; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2927; B =3202; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6101; B =7618; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7898; B =5737; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8390; B =2606; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6700; B =1502; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8481; B =7415; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2095; B =2106; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8266; B =1731; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9736; B =7160; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5113; B =9154; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8466; B =3805; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6175; B =4119; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1581; B =3961; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4708; B =3363; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7611; B =5901; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0293; B =5356; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3547; B =3889; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0695; B =0367; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5336; B =9836; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5988; B =5223; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6637; B =0340; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1443; B =2993; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9130; B =1602; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3467; B =8436; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9554; B =5561; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0387; B =1261; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2931; B =2617; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6222; B =5757; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4279; B =1060; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9840; B =5622; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3162; B =4383; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2538; B =8306; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7495; B =9518; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7603; B =3599; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8490; B =6870; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7463; B =5822; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9427; B =9893; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7618; B =6422; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5546; B =7591; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0485; B =7323; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6238; B =1901; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4703; B =7240; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2131; B =2011; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5038; B =0721; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6272; B =4206; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2562; B =4565; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9289; B =8656; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4244; B =0868; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9322; B =2919; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1449; B =5997; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3678; B =7046; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9897; B =2938; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8971; B =1715; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2320; B =2183; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5436; B =7727; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1502; B =7086; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4323; B =3527; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9845; B =8120; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0879; B =1503; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5498; B =6371; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4442; B =2095; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3073; B =1971; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9281; B =0823; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7771; B =3032; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2056; B =2152; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1684; B =9550; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4549; B =7761; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9541; B =7771; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0074; B =4949; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1153; B =0117; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8174; B =8175; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2894; B =1702; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2691; B =9660; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2753; B =5546; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8458; B =5837; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1844; B =8122; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9959; B =3081; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9655; B =7637; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7764; B =4513; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9798; B =9225; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9771; B =4259; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5019; B =1277; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4797; B =4529; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9291; B =2171; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9502; B =3879; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2735; B =7225; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0396; B =3796; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2621; B =5481; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0292; B =9601; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0708; B =4207; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0970; B =0666; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8647; B =1825; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0487; B =4299; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5150; B =2233; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5787; B =5362; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5712; B =9154; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6745; B =9735; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2962; B =3415; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5179; B =8876; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3689; B =0233; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0618; B =0156; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5598; B =8531; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6246; B =6407; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6287; B =1390; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9731; B =7852; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7966; B =5747; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4056; B =2336; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3193; B =6817; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9285; B =7097; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5214; B =0582; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7304; B =0436; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9775; B =8734; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4637; B =4798; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6703; B =3721; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5212; B =3312; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2285; B =3554; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7505; B =0565; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9782; B =7020; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5357; B =1624; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4479; B =6956; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2601; B =3736; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8470; B =0632; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3044; B =5514; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0010; B =6895; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9878; B =0755; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2656; B =6748; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5777; B =2489; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6421; B =9553; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5367; B =4949; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7768; B =2491; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4850; B =7654; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1412; B =2411; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6275; B =3792; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7389; B =1598; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8862; B =8129; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1163; B =4103; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5009; B =7304; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7907; B =4708; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1430; B =7582; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1423; B =3273; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2655; B =6210; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =3501; B =8944; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =6396; B =4928; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9106; B =8198; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2921; B =8876; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4270; B =9848; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4907; B =0061; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1343; B =5845; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8668; B =1811; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7955; B =9979; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7927; B =6495; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2289; B =9455; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =9906; B =6717; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =8061; B =2487; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =0004; B =7132; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7125; B =9271; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =7770; B =1760; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =1061; B =3452; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =5672; B =9107; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =2681; B =7942; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100 A =4540; B =6706; Sub = 1;Op1 = 1; Op2 = 1; Cin = 0; Less = 0;
			#100
			
			$display($time, ,"A=%d, B=%d, Cin=%b, F=%d, Cout=%b, Set=%b, Sub=%b, Op1=%b, Op2=%b, Less=%b", A, B, Cin,F, Cout, Set, Sub, Op1, Op2, Less);
		end
endmodule


module ALU16(F, Cout, Set, Less, A, B, Cin, Sub, Op1, Op2);//code for 16, 1-bit ALUs wired together

	output [15:0] F, Cout, Set;
	input [15:0] A, B;
	input Op1, Op2, Sub, Cin, Less;

	return r0 (F[0], Cout[0], Set[0], Set[15], A[0], B[0], Sub, Sub, Op1, Op2);
	return r1 (F[1], Cout[1], Set[1], 0, A[1], B[1], Cout[0], Sub, Op1, Op2);
	return r2 (F[2], Cout[2], Set[2], 0, A[2], B[2], Cout[1], Sub, Op1, Op2);
	return r3 (F[3], Cout[3], Set[3], 0, A[3], B[3], Cout[2], Sub, Op1, Op2);
	return r4 (F[4], Cout[4], Set[4], 0, A[4], B[4], Cout[3], Sub, Op1, Op2);
	return r5 (F[5], Cout[5], Set[5], 0, A[5], B[5], Cout[4], Sub, Op1, Op2);
	return r6 (F[6], Cout[6], Set[6], 0, A[6], B[6], Cout[5], Sub, Op1, Op2);
	return r7 (F[7], Cout[7], Set[7], 0, A[7], B[7], Cout[6], Sub, Op1, Op2);
	return r8 (F[8], Cout[8], Set[8], 0, A[8], B[8], Cout[7], Sub, Op1, Op2);
	return r9 (F[9], Cout[9], Set[9], 0, A[9], B[9], Cout[8], Sub, Op1, Op2);
	return r10 (F[10], Cout[10], Set[10], 0, A[10], B[10], Cout[9], Sub, Op1, Op2);
	return r11 (F[11], Cout[11], Set[11], 0, A[11], B[11], Cout[10], Sub, Op1, Op2);
	return r12 (F[12], Cout[12], Set[12], 0, A[12], B[12], Cout[11], Sub, Op1, Op2);
	return r13 (F[13], Cout[13], Set[13], 0, A[13], B[13], Cout[12], Sub, Op1, Op2);
	return r14 (F[14], Cout[14], Set[14], 0, A[14], B[14], Cout[13], Sub, Op1, Op2);
	return r15 (F[15], Cout[15], Set[15], 0, A[15], B[15], Cout[14], Sub, Op1, Op2);

endmodule

module return(F,Cout,Set,Less,A,B,Cin,Sub,Op1,Op2);//Code for a 1-bit ALU

   output F,Cout, Set;
   input  A, B, Cin, Sub, Op1, Op2, Less;
   wire   w1, w2, w3, w4;
 
   fulladder FA (Set, Cout, A, w4, Cin);
   four_to_one_mux F1 (F, w1, w2, Set, Less, Op1, Op2);
   xor #1 G4(w4, Sub, B);
   and #1 G1(w1, A, B);
   or #1 G2(w2, A, B);
 
endmodule


module four_to_one_mux(F, A, B, C, D, S1, S2); //code for a basic 4-1 mux used in a 1-bit ALU
	
	wire w1, w2, w3, w4, w5, w6;
	input A, B, C, D, S1, S2;
	output F;
	
	not #1 G1(w1, S1);
	not #1 G2(w2, S2);
	and #1 G3(w3, A, w1, w2);
	and #1 G4(w4, B, S2, w1);
	and #1 G5(w5, C, S1, w2);
	and #1 G6(w6, D, S1, S2);
	or #1 G7(F, w3, w4, w5, w6);

endmodule

module fulladder(S,Cout,A,B,Cin);//code for a full adder with a 1 nanosecond delay

	output S, Cout;
	input A, B, Cin;
	wire w1, w2, w3, w4, w5;

	xor #1 G1(w1, A, B);
	xor #1 G6(S, w1, Cin);
	and #1 G2(w2, A, Cin);
	and #1 G3(w3, B, Cin);
	and #1 G4(w4, A, B);
	or #1 G5(Cout, w2, w3, w4);
endmodule